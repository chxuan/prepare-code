module moduleName (
    ports
);
    
endmodule